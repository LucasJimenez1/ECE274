`timescale 1ns / 1ps
module Lab5_top_level(Clk, Rst, go, done, sum);
    input Clk; //clock
    input Rst; //reset
    input go;
    output done;
    output sum;

endmodule
